module ALU (clk, rst, Op_code, Addr_1, Addr_2, Output);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [31:0] Op_code;
  input  wire [31:0] Addr_1;
  input  wire [31:0] Addr_2;
  output  wire [15:0] Output;

  TC_Add # (.UUID(64'd771736472665924867 ^ UUID), .BIT_WIDTH(64'd32)) Add32_0 (.in0(wire_12), .in1(wire_5), .ci(1'd0), .out(wire_35), .co());
  TC_Switch # (.UUID(64'd4291707569989912967 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_1 (.en(wire_19), .in(wire_35), .out(wire_4_10));
  TC_And # (.UUID(64'd2367903160720416068 ^ UUID), .BIT_WIDTH(64'd64)) And64_2 (.in0({{32{1'b0}}, wire_23 }), .in1({{32{1'b0}}, wire_33 }), .out(wire_1));
  TC_Constant # (.UUID(64'd3702637439539675981 ^ UUID), .BIT_WIDTH(64'd32), .value(32'hFF)) Constant32_3 (.out(wire_33));
  TC_Equal # (.UUID(64'd3307467026970206130 ^ UUID), .BIT_WIDTH(64'd32)) Equal32_4 (.in0(wire_1[31:0]), .in1(wire_31), .out(wire_19));
  TC_Constant # (.UUID(64'd2969093834876989049 ^ UUID), .BIT_WIDTH(64'd32), .value(32'h0)) Constant32_5 (.out(wire_31));
  TC_Add # (.UUID(64'd1192413511963083168 ^ UUID), .BIT_WIDTH(64'd32)) Add32_6 (.in0(wire_12), .in1(wire_17), .ci(1'd0), .out(wire_20), .co());
  TC_Switch # (.UUID(64'd3466348840251439509 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_7 (.en(wire_28), .in(wire_20), .out(wire_4_9));
  TC_Equal # (.UUID(64'd982387346584071466 ^ UUID), .BIT_WIDTH(64'd32)) Equal32_8 (.in0(wire_1[31:0]), .in1(wire_29), .out(wire_28));
  TC_Constant # (.UUID(64'd4281366940539241251 ^ UUID), .BIT_WIDTH(64'd32), .value(32'h1)) Constant32_9 (.out(wire_29));
  TC_Neg # (.UUID(64'd2104763954609761425 ^ UUID), .BIT_WIDTH(64'd32)) Neg32_10 (.in(wire_5), .out(wire_17));
  TC_Switch # (.UUID(64'd454292827248976047 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_11 (.en(wire_15), .in(wire_2), .out(wire_4_8));
  TC_Equal # (.UUID(64'd1886273917479343232 ^ UUID), .BIT_WIDTH(64'd32)) Equal32_12 (.in0(wire_1[31:0]), .in1(wire_3), .out(wire_15));
  TC_Constant # (.UUID(64'd1036248000938172543 ^ UUID), .BIT_WIDTH(64'd32), .value(32'h2)) Constant32_13 (.out(wire_3));
  TC_And # (.UUID(64'd2966261516107634040 ^ UUID), .BIT_WIDTH(64'd32)) And32_14 (.in0(wire_12), .in1(wire_5), .out(wire_2));
  TC_Switch # (.UUID(64'd4244556451358743428 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_15 (.en(wire_16), .in(wire_32), .out(wire_4_7));
  TC_Equal # (.UUID(64'd2378019975791647168 ^ UUID), .BIT_WIDTH(64'd32)) Equal32_16 (.in0(wire_1[31:0]), .in1(wire_8), .out(wire_16));
  TC_Constant # (.UUID(64'd3649162839773976333 ^ UUID), .BIT_WIDTH(64'd32), .value(32'h3)) Constant32_17 (.out(wire_8));
  TC_Or # (.UUID(64'd1919012726298350117 ^ UUID), .BIT_WIDTH(64'd32)) Or32_18 (.in0(wire_12), .in1(wire_5), .out(wire_32));
  TC_Switch # (.UUID(64'd279021741894509172 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_19 (.en(wire_37), .in(wire_18), .out(wire_4_6));
  TC_Equal # (.UUID(64'd2683582231972257440 ^ UUID), .BIT_WIDTH(64'd32)) Equal32_20 (.in0(wire_1[31:0]), .in1(wire_10), .out(wire_37));
  TC_Constant # (.UUID(64'd2598932003380171208 ^ UUID), .BIT_WIDTH(64'd32), .value(32'h4)) Constant32_21 (.out(wire_10));
  TC_Nand # (.UUID(64'd4271646140554606194 ^ UUID), .BIT_WIDTH(64'd32)) Nand32_22 (.in0(wire_12), .in1(wire_5), .out(wire_18));
  TC_Switch # (.UUID(64'd4105564870275111942 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_23 (.en(wire_26), .in(wire_21), .out(wire_4_5));
  TC_Equal # (.UUID(64'd3962148131258842660 ^ UUID), .BIT_WIDTH(64'd32)) Equal32_24 (.in0(wire_1[31:0]), .in1(wire_39), .out(wire_26));
  TC_Constant # (.UUID(64'd3292953784274058964 ^ UUID), .BIT_WIDTH(64'd32), .value(32'h5)) Constant32_25 (.out(wire_39));
  TC_Nor # (.UUID(64'd2094435172533730788 ^ UUID), .BIT_WIDTH(64'd32)) Nor32_26 (.in0(wire_12), .in1(wire_5), .out(wire_21));
  TC_Switch # (.UUID(64'd4395527959694623491 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_27 (.en(wire_14), .in(wire_11), .out(wire_4_4));
  TC_Equal # (.UUID(64'd2728722859468860567 ^ UUID), .BIT_WIDTH(64'd32)) Equal32_28 (.in0(wire_1[31:0]), .in1(wire_27), .out(wire_14));
  TC_Constant # (.UUID(64'd2814141242211950990 ^ UUID), .BIT_WIDTH(64'd32), .value(32'h6)) Constant32_29 (.out(wire_27));
  TC_Xor # (.UUID(64'd1561626617431980233 ^ UUID), .BIT_WIDTH(64'd32)) Xor32_30 (.in0(wire_12), .in1(wire_5), .out(wire_11));
  TC_Switch # (.UUID(64'd25380029634364728 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_31 (.en(wire_9), .in(wire_36), .out(wire_4_3));
  TC_Equal # (.UUID(64'd1804665057419404565 ^ UUID), .BIT_WIDTH(64'd32)) Equal32_32 (.in0(wire_1[31:0]), .in1(wire_22), .out(wire_9));
  TC_Constant # (.UUID(64'd1036449072606840649 ^ UUID), .BIT_WIDTH(64'd32), .value(32'h7)) Constant32_33 (.out(wire_22));
  TC_Switch # (.UUID(64'd1731737387117890663 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_34 (.en(wire_30), .in(wire_7), .out(wire_4_1));
  TC_Equal # (.UUID(64'd3023334011462849504 ^ UUID), .BIT_WIDTH(64'd32)) Equal32_35 (.in0(wire_1[31:0]), .in1(wire_0), .out(wire_30));
  TC_Constant # (.UUID(64'd1980186390380277652 ^ UUID), .BIT_WIDTH(64'd32), .value(32'h8)) Constant32_36 (.out(wire_0));
  TC_Shl # (.UUID(64'd354489379800897438 ^ UUID), .BIT_WIDTH(64'd32)) Shl32_37 (.in(wire_12), .shift(wire_5[7:0]), .out(wire_36));
  TC_Switch # (.UUID(64'd2738600531205630654 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_38 (.en(wire_38), .in(wire_13), .out(wire_4_0));
  TC_Equal # (.UUID(64'd3712194815650869653 ^ UUID), .BIT_WIDTH(64'd32)) Equal32_39 (.in0(wire_1[31:0]), .in1(wire_6), .out(wire_38));
  TC_Constant # (.UUID(64'd1535763231293589767 ^ UUID), .BIT_WIDTH(64'd32), .value(32'h9)) Constant32_40 (.out(wire_6));
  TC_Shr # (.UUID(64'd4428106322157092189 ^ UUID), .BIT_WIDTH(64'd32)) Shr32_41 (.in(wire_12), .shift(wire_5[7:0]), .out(wire_7));
  TC_Switch # (.UUID(64'd2602867552618789742 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_42 (.en(wire_24), .in(wire_34), .out(wire_4_2));
  TC_Equal # (.UUID(64'd833107010798282109 ^ UUID), .BIT_WIDTH(64'd32)) Equal32_43 (.in0(wire_1[31:0]), .in1(wire_25), .out(wire_24));
  TC_Constant # (.UUID(64'd2748849295724651539 ^ UUID), .BIT_WIDTH(64'd32), .value(32'hA)) Constant32_44 (.out(wire_25));
  TC_Not # (.UUID(64'd662502363542981586 ^ UUID), .BIT_WIDTH(64'd32)) Not32_45 (.in(wire_12), .out(wire_13));
  TC_Neg # (.UUID(64'd1903017984973985502 ^ UUID), .BIT_WIDTH(64'd32)) Neg32_46 (.in(wire_12), .out(wire_34));

  wire [31:0] wire_0;
  wire [63:0] wire_1;
  wire [31:0] wire_2;
  wire [31:0] wire_3;
  wire [31:0] wire_4;
  wire [31:0] wire_4_0;
  wire [31:0] wire_4_1;
  wire [31:0] wire_4_2;
  wire [31:0] wire_4_3;
  wire [31:0] wire_4_4;
  wire [31:0] wire_4_5;
  wire [31:0] wire_4_6;
  wire [31:0] wire_4_7;
  wire [31:0] wire_4_8;
  wire [31:0] wire_4_9;
  wire [31:0] wire_4_10;
  assign wire_4 = wire_4_0|wire_4_1|wire_4_2|wire_4_3|wire_4_4|wire_4_5|wire_4_6|wire_4_7|wire_4_8|wire_4_9|wire_4_10;
  assign Output = wire_4[15:0];
  wire [31:0] wire_5;
  assign wire_5 = Addr_2;
  wire [31:0] wire_6;
  wire [31:0] wire_7;
  wire [31:0] wire_8;
  wire [0:0] wire_9;
  wire [31:0] wire_10;
  wire [31:0] wire_11;
  wire [31:0] wire_12;
  assign wire_12 = Addr_1;
  wire [31:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [0:0] wire_16;
  wire [31:0] wire_17;
  wire [31:0] wire_18;
  wire [0:0] wire_19;
  wire [31:0] wire_20;
  wire [31:0] wire_21;
  wire [31:0] wire_22;
  wire [31:0] wire_23;
  assign wire_23 = Op_code;
  wire [0:0] wire_24;
  wire [31:0] wire_25;
  wire [0:0] wire_26;
  wire [31:0] wire_27;
  wire [0:0] wire_28;
  wire [31:0] wire_29;
  wire [0:0] wire_30;
  wire [31:0] wire_31;
  wire [31:0] wire_32;
  wire [31:0] wire_33;
  wire [31:0] wire_34;
  wire [31:0] wire_35;
  wire [31:0] wire_36;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  wire [31:0] wire_39;

endmodule
